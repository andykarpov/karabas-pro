-- megafunction wizard: %ALTCLKCTRL%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altclkctrl 

-- ============================================================
-- File Name: clk_ctrl2.vhd
-- Megafunction Name(s):
-- 			altclkctrl
--
-- Simulation Library Files(s):
-- 			cycloneive
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 13.0.1 Build 232 06/12/2013 SP 1 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2013 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


--altclkctrl CBX_AUTO_BLACKBOX="ALL" CLOCK_TYPE="Global Clock" DEVICE_FAMILY="Cyclone IV E" ENA_REGISTER_MODE="falling edge" USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION="ON" clkselect ena inclk outclk
--VERSION_BEGIN 13.0 cbx_altclkbuf 2013:06:12:18:03:43:SJ cbx_cycloneii 2013:06:12:18:03:43:SJ cbx_lpm_add_sub 2013:06:12:18:03:43:SJ cbx_lpm_compare 2013:06:12:18:03:43:SJ cbx_lpm_decode 2013:06:12:18:03:43:SJ cbx_lpm_mux 2013:06:12:18:03:43:SJ cbx_mgl 2013:06:12:18:05:10:SJ cbx_stratix 2013:06:12:18:03:43:SJ cbx_stratixii 2013:06:12:18:03:43:SJ cbx_stratixiii 2013:06:12:18:03:43:SJ cbx_stratixv 2013:06:12:18:03:43:SJ  VERSION_END

 LIBRARY cycloneive;
 USE cycloneive.all;

--synthesis_resources = clkctrl 1 reg 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  clk_ctrl2_altclkctrl_9gi IS 
	 PORT 
	 ( 
		 clkselect	:	IN  STD_LOGIC_VECTOR (1 DOWNTO 0) := (OTHERS => '0');
		 ena	:	IN  STD_LOGIC := '1';
		 inclk	:	IN  STD_LOGIC_VECTOR (3 DOWNTO 0) := (OTHERS => '0');
		 outclk	:	OUT  STD_LOGIC
	 ); 
 END clk_ctrl2_altclkctrl_9gi;

 ARCHITECTURE RTL OF clk_ctrl2_altclkctrl_9gi IS

	 ATTRIBUTE synthesis_clearbox : natural;
	 ATTRIBUTE synthesis_clearbox OF RTL : ARCHITECTURE IS 2;
	 ATTRIBUTE ALTERA_ATTRIBUTE : string;
	 SIGNAL	 ena_reg	:	STD_LOGIC
	 -- synopsys translate_off
	  := '1'
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF ena_reg : SIGNAL IS "POWER_UP_LEVEL=HIGH";

	 SIGNAL  wire_ena_reg_w_lg_q6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 select_reg	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 ATTRIBUTE ALTERA_ATTRIBUTE OF select_reg : SIGNAL IS "POWER_UP_LEVEL=LOW";

	 SIGNAL  wire_select_reg_w_q_range12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_select_reg_w_q_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_clkctrl1_w_lg_outclk5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_clkctrl1_clkselect	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_clkctrl1_outclk	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_select_enable_wire_range14w20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_clkselect_wire_range13w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_clkselect_wire_range18w19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  clkselect_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  inclk_wire :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  select_enable_wire :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_clkselect_wire_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_clkselect_wire_range3w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_w_clkselect_wire_range18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_select_enable_wire_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  cycloneive_clkctrl
	 GENERIC 
	 (
		clock_type	:	STRING;
		ena_register_mode	:	STRING := "falling edge";
		lpm_type	:	STRING := "cycloneive_clkctrl"
	 );
	 PORT
	 ( 
		clkselect	:	IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		ena	:	IN STD_LOGIC;
		inclk	:	IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		outclk	:	OUT STD_LOGIC
	 ); 
	 END COMPONENT;
 BEGIN

	wire_vcc <= '1';
	wire_w_lg_w_select_enable_wire_range14w20w(0) <= wire_w_select_enable_wire_range14w(0) OR wire_w_lg_w_clkselect_wire_range18w19w(0);
	wire_w_lg_w_clkselect_wire_range13w15w(0) <= wire_w_clkselect_wire_range13w(0) XOR wire_select_reg_w_q_range12w(0);
	wire_w_lg_w_clkselect_wire_range18w19w(0) <= wire_w_clkselect_wire_range18w(0) XOR wire_select_reg_w_q_range17w(0);
	clkselect_wire <= ( clkselect);
	inclk_wire <= ( inclk);
	outclk <= (wire_clkctrl1_outclk AND ena_reg);
	select_enable_wire <= ( wire_w_lg_w_select_enable_wire_range14w20w & wire_w_lg_w_clkselect_wire_range13w15w);
	wire_w_clkselect_wire_range13w(0) <= clkselect_wire(0);
	wire_w_clkselect_wire_range3w <= clkselect_wire(1 DOWNTO 0);
	wire_w_clkselect_wire_range18w(0) <= clkselect_wire(1);
	wire_w_select_enable_wire_range14w(0) <= select_enable_wire(0);
	PROCESS (wire_clkctrl1_outclk)
	BEGIN
		IF (wire_clkctrl1_outclk = '0' AND wire_clkctrl1_outclk'event) THEN ena_reg <= (ena AND (NOT select_enable_wire(1)));
		END IF;
	END PROCESS;
	PROCESS (wire_clkctrl1_outclk)
	BEGIN
		IF (wire_clkctrl1_outclk = '0' AND wire_clkctrl1_outclk'event) THEN 
			IF (ena_reg = '0') THEN select_reg <= wire_w_clkselect_wire_range3w;
			END IF;
		END IF;
	END PROCESS;
	wire_select_reg_w_q_range12w(0) <= select_reg(0);
	wire_select_reg_w_q_range17w(0) <= select_reg(1);
	wire_clkctrl1_w_lg_outclk5w(0) <= NOT wire_clkctrl1_outclk;
	wire_clkctrl1_clkselect <= ( select_reg);
	clkctrl1 :  cycloneive_clkctrl
	  GENERIC MAP (
		clock_type => "Global Clock"
	  )
	  PORT MAP ( 
		clkselect => wire_clkctrl1_clkselect,
		ena => wire_vcc,
		inclk => inclk_wire,
		outclk => wire_clkctrl1_outclk
	  );

 END RTL; --clk_ctrl2_altclkctrl_9gi
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY clk_ctrl2 IS
	PORT
	(
		clkselect		: IN STD_LOGIC  := '0';
		inclk0x		: IN STD_LOGIC ;
		inclk1x		: IN STD_LOGIC ;
		outclk		: OUT STD_LOGIC 
	);
END clk_ctrl2;


ARCHITECTURE RTL OF clk_ctrl2 IS

	ATTRIBUTE synthesis_clearbox: natural;
	ATTRIBUTE synthesis_clearbox OF RTL: ARCHITECTURE IS 2;
	ATTRIBUTE clearbox_macroname: string;
	ATTRIBUTE clearbox_macroname OF RTL: ARCHITECTURE IS "altclkctrl";
	ATTRIBUTE clearbox_defparam: string;
	ATTRIBUTE clearbox_defparam OF RTL: ARCHITECTURE IS "ena_register_mode=falling edge;intended_device_family=Cyclone IV E;use_glitch_free_switch_over_implementation=ON;clock_type=Global Clock;";
	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC ;
	SIGNAL sub_wire2	: STD_LOGIC_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire3_bv	: BIT_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (0 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC ;
	SIGNAL sub_wire5	: STD_LOGIC ;
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (3 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC ;
	SIGNAL sub_wire8_bv	: BIT_VECTOR (1 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (1 DOWNTO 0);



	COMPONENT clk_ctrl2_altclkctrl_9gi
	PORT (
			clkselect	: IN STD_LOGIC_VECTOR (1 DOWNTO 0);
			ena	: IN STD_LOGIC ;
			inclk	: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
			outclk	: OUT STD_LOGIC 
	);
	END COMPONENT;

BEGIN
	sub_wire3_bv(0 DOWNTO 0) <= "0";
	sub_wire3    <= To_stdlogicvector(sub_wire3_bv);
	sub_wire4    <= '1';
	sub_wire8_bv(1 DOWNTO 0) <= "00";
	sub_wire8    <= To_stdlogicvector(sub_wire8_bv);
	sub_wire7    <= inclk1x;
	outclk    <= sub_wire0;
	sub_wire1    <= clkselect;
	sub_wire2    <= sub_wire3(0 DOWNTO 0) & sub_wire1;
	sub_wire5    <= inclk0x;
	sub_wire6    <= sub_wire8(1 DOWNTO 0) & sub_wire7 & sub_wire5;

	clk_ctrl2_altclkctrl_9gi_component : clk_ctrl2_altclkctrl_9gi
	PORT MAP (
		clkselect => sub_wire2,
		ena => sub_wire4,
		inclk => sub_wire6,
		outclk => sub_wire0
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: PRIVATE: clock_inputs NUMERIC "2"
-- Retrieval info: CONSTANT: ENA_REGISTER_MODE STRING "falling edge"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: USE_GLITCH_FREE_SWITCH_OVER_IMPLEMENTATION STRING "ON"
-- Retrieval info: CONSTANT: clock_type STRING "Global Clock"
-- Retrieval info: USED_PORT: clkselect 0 0 0 0 INPUT GND "clkselect"
-- Retrieval info: USED_PORT: inclk0x 0 0 0 0 INPUT NODEFVAL "inclk0x"
-- Retrieval info: USED_PORT: inclk1x 0 0 0 0 INPUT NODEFVAL "inclk1x"
-- Retrieval info: USED_PORT: outclk 0 0 0 0 OUTPUT NODEFVAL "outclk"
-- Retrieval info: CONNECT: @clkselect 0 0 1 1 GND 0 0 0 0
-- Retrieval info: CONNECT: @clkselect 0 0 1 0 clkselect 0 0 0 0
-- Retrieval info: CONNECT: @ena 0 0 0 0 VCC 0 0 0 0
-- Retrieval info: CONNECT: @inclk 0 0 2 2 GND 0 0 2 0
-- Retrieval info: CONNECT: @inclk 0 0 1 0 inclk0x 0 0 0 0
-- Retrieval info: CONNECT: @inclk 0 0 1 1 inclk1x 0 0 0 0
-- Retrieval info: CONNECT: outclk 0 0 0 0 @outclk 0 0 0 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL clk_ctrl2.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL clk_ctrl2.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL clk_ctrl2.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL clk_ctrl2.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL clk_ctrl2_inst.vhd FALSE
-- Retrieval info: LIB_FILE: cycloneive
