//----------------------------------------------------------------------------
//  A-Z80 CPU Copyright (C) 2014,2017  Goran Devic, www.baltazarstudios.com
//
//  This program is free software; you can redistribute it and/or modify it
//  under the terms of the GNU General Public License as published by the Free
//  Software Foundation; either version 2 of the License, or (at your option)
//  any later version.
//
//  This program is distributed in the hope that it will be useful, but WITHOUT
//  ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or
//  FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License for
//  more details.
//----------------------------------------------------------------------------
// Automatically generated by gencompile.py

reg ctl_reg_gp_sel_pla17npla50M1T1_2;
reg ctl_reg_gp_hilo_pla17npla50M1T1_3;
reg ctl_reg_sys_hilo_pla17npla50M2T1_3;
reg ctl_reg_sys_hilo_pla17npla50M2T2_4;
reg ctl_reg_gp_sel_pla61npla58npla59M1T1_2;
reg ctl_reg_gp_hilo_pla61npla58npla59M1T1_3;
reg ctl_reg_gp_sel_pla61npla58npla59M1T4_3;
reg ctl_reg_gp_hilo_pla61npla58npla59M1T4_4;
reg ctl_reg_gp_sel_use_ixiypla58M1T1_2;
reg ctl_reg_gp_hilo_use_ixiypla58M1T1_3;
reg ctl_reg_sys_hilo_use_ixiypla58M2T1_3;
reg ctl_reg_sys_hilo_use_ixiypla58M2T2_4;
reg ctl_reg_gp_sel_nuse_ixiypla58M1T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla58M1T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla58M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla58M2T1_3;
reg ctl_reg_sys_hilo_use_ixiypla59M2T1_3;
reg ctl_reg_sys_hilo_use_ixiypla59M2T2_4;
reg ctl_reg_gp_sel_nuse_ixiypla59M1T4_4;
reg ctl_reg_gp_hilo_nuse_ixiypla59M1T4_5;
reg ctl_reg_gp_sel_nuse_ixiypla59M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla59M2T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla59M4T1_3;
reg ctl_reg_gp_hilo_nuse_ixiypla59M4T1_4;
reg ctl_reg_sys_hilo_pla40M2T1_3;
reg ctl_reg_sys_hilo_pla40M2T2_4;
reg ctl_reg_sys_hilo_pla40M3T1_3;
reg ctl_reg_sys_hilo_pla40M3T2_4;
reg ctl_reg_sys_hilo_pla50npla40M2T1_3;
reg ctl_reg_sys_hilo_pla50npla40M2T2_4;
reg ctl_reg_gp_sel_pla50npla40M3T1_2;
reg ctl_reg_gp_hilo_pla50npla40M3T1_3;
reg ctl_reg_gp_sel_pla8pla13M1T4_4;
reg ctl_reg_gp_hilo_pla8pla13M1T4_5;
reg ctl_reg_gp_sel_pla8pla13M2T1_2;
reg ctl_reg_gp_hilo_pla8pla13M2T1_3;
reg ctl_reg_sys_hilo_pla8pla13M2T2_4;
reg ctl_reg_gp_sel_pla8npla13M1T1_2;
reg ctl_reg_gp_hilo_pla8npla13M1T1_3;
reg ctl_reg_gp_sel_pla8npla13M2T1_2;
reg ctl_reg_gp_hilo_pla8npla13M2T1_3;
reg ctl_reg_sys_hilo_pla8npla13M2T2_4;
reg ctl_reg_sys_hilo_pla38pla13M2T1_3;
reg ctl_reg_sys_hilo_pla38pla13M2T2_4;
reg ctl_reg_sys_hilo_pla38pla13M2T3_6;
reg ctl_reg_sys_hilo_pla38pla13M3T1_3;
reg ctl_reg_sys_hilo_pla38pla13M3T2_4;
reg ctl_reg_sys_hilo_pla38pla13M3T3_5;
reg ctl_reg_sys_hilo_pla38pla13M3T3_10;
reg ctl_reg_gp_sel_pla38pla13M4T1_3;
reg ctl_reg_gp_hilo_pla38pla13M4T1_4;
reg ctl_reg_sys_hilo_pla38pla13M4T2_4;
reg ctl_reg_gp_sel_pla38npla13M1T1_2;
reg ctl_reg_gp_hilo_pla38npla13M1T1_3;
reg ctl_reg_sys_hilo_pla38npla13M2T1_3;
reg ctl_reg_sys_hilo_pla38npla13M2T2_4;
reg ctl_reg_sys_hilo_pla38npla13M2T3_6;
reg ctl_reg_sys_hilo_pla38npla13M3T1_3;
reg ctl_reg_sys_hilo_pla38npla13M3T2_4;
reg ctl_reg_sys_hilo_pla38npla13M3T3_6;
reg ctl_reg_sys_hilo_pla38npla13M4T1_3;
reg ctl_reg_sys_hilo_pla38npla13M4T2_4;
reg ctl_reg_gp_sel_pla83M1T1_2;
reg ctl_reg_gp_hilo_pla83M1T1_3;
reg ctl_pf_sel_pla83M1T1_19;
reg ctl_reg_gp_sel_pla83M1T2_2;
reg ctl_reg_gp_hilo_pla83M1T2_3;
reg ctl_reg_gp_sel_pla83M1T3_1;
reg ctl_reg_gp_hilo_pla83M1T3_2;
reg ctl_reg_sys_hilo_pla83M1T4_3;
reg ctl_reg_gp_sel_pla57M1T3_1;
reg ctl_reg_gp_hilo_pla57M1T3_2;
reg ctl_reg_sys_hilo_pla57M1T4_4;
reg ctl_reg_gp_sel_pla7M1T1_2;
reg ctl_reg_gp_hilo_pla7M1T1_3;
reg ctl_reg_sys_hilo_pla7M2T1_3;
reg ctl_reg_sys_hilo_pla7M2T2_4;
reg ctl_reg_sys_hilo_pla7M3T1_3;
reg ctl_reg_gp_sel_pla7M3T1_6;
reg ctl_reg_gp_hilo_pla7M3T1_7;
reg ctl_reg_sys_hilo_pla7M3T2_4;
reg ctl_reg_sys_hilo_pla30pla13M2T1_3;
reg ctl_reg_sys_hilo_pla30pla13M2T2_4;
reg ctl_reg_sys_hilo_pla30pla13M2T3_6;
reg ctl_reg_sys_hilo_pla30pla13M3T1_3;
reg ctl_reg_sys_hilo_pla30pla13M3T2_4;
reg ctl_reg_sys_hilo_pla30pla13M3T3_5;
reg ctl_reg_sys_hilo_pla30pla13M3T3_10;
reg ctl_reg_gp_sel_pla30pla13M4T1_3;
reg ctl_reg_gp_hilo_pla30pla13M4T1_4;
reg ctl_reg_sys_hilo_pla30pla13M4T2_4;
reg ctl_reg_sys_hilo_pla30pla13M4T3_5;
reg ctl_reg_gp_sel_pla30pla13M5T1_3;
reg ctl_reg_gp_hilo_pla30pla13M5T1_4;
reg ctl_reg_sys_hilo_pla30pla13M5T2_4;
reg ctl_reg_sys_hilo_pla30npla13M2T1_3;
reg ctl_reg_sys_hilo_pla30npla13M2T2_4;
reg ctl_reg_sys_hilo_pla30npla13M2T3_6;
reg ctl_reg_sys_hilo_pla30npla13M3T1_3;
reg ctl_reg_sys_hilo_pla30npla13M3T2_4;
reg ctl_reg_sys_hilo_pla30npla13M3T3_6;
reg ctl_reg_sys_hilo_pla30npla13M4T1_3;
reg ctl_reg_sys_hilo_pla30npla13M4T2_4;
reg ctl_reg_gp_sel_pla30npla13M4T3_5;
reg ctl_reg_gp_hilo_pla30npla13M4T3_6;
reg ctl_reg_sys_hilo_pla30npla13M5T1_3;
reg ctl_reg_sys_hilo_pla30npla13M5T2_4;
reg ctl_reg_gp_sel_pla30npla13M5T3_4;
reg ctl_reg_gp_hilo_pla30npla13M5T3_5;
reg ctl_reg_sys_hilo_pla31pla33M2T1_3;
reg ctl_reg_sys_hilo_pla31pla33M2T2_4;
reg ctl_reg_sys_hilo_pla31pla33M2T3_6;
reg ctl_reg_sys_hilo_pla31pla33M3T1_3;
reg ctl_reg_sys_hilo_pla31pla33M3T2_4;
reg ctl_reg_sys_hilo_pla31pla33M3T3_5;
reg ctl_reg_sys_hilo_pla31pla33M3T3_10;
reg ctl_reg_gp_sel_pla31pla33M4T1_3;
reg ctl_reg_gp_hilo_pla31pla33M4T1_4;
reg ctl_reg_sys_hilo_pla31pla33M4T2_4;
reg ctl_reg_sys_hilo_pla31pla33M4T3_5;
reg ctl_reg_gp_sel_pla31pla33M5T1_3;
reg ctl_reg_gp_hilo_pla31pla33M5T1_4;
reg ctl_reg_sys_hilo_pla31pla33M5T2_4;
reg ctl_reg_sys_hilo_pla31npla33M2T1_3;
reg ctl_reg_sys_hilo_pla31npla33M2T2_4;
reg ctl_reg_sys_hilo_pla31npla33M2T3_6;
reg ctl_reg_sys_hilo_pla31npla33M3T1_3;
reg ctl_reg_sys_hilo_pla31npla33M3T2_4;
reg ctl_reg_sys_hilo_pla31npla33M3T3_6;
reg ctl_reg_sys_hilo_pla31npla33M4T1_3;
reg ctl_reg_sys_hilo_pla31npla33M4T2_4;
reg ctl_reg_gp_sel_pla31npla33M4T3_5;
reg ctl_reg_gp_hilo_pla31npla33M4T3_6;
reg ctl_reg_sys_hilo_pla31npla33M5T1_3;
reg ctl_reg_sys_hilo_pla31npla33M5T2_4;
reg ctl_reg_gp_sel_pla31npla33M5T3_4;
reg ctl_reg_gp_hilo_pla31npla33M5T3_5;
reg ctl_reg_gp_sel_pla5M1T4_2;
reg ctl_reg_gp_hilo_pla5M1T4_3;
reg ctl_reg_gp_sel_pla5M1T5_2;
reg ctl_reg_gp_hilo_pla5M1T5_3;
reg ctl_reg_gp_sel_pla23pla16M1T5_4;
reg ctl_reg_gp_hilo_pla23pla16M1T5_5;
reg ctl_reg_gp_sel_pla23pla16M2T1_5;
reg ctl_reg_gp_hilo_pla23pla16M2T1_6;
reg ctl_reg_gp_sel_pla23pla16M2T2_3;
reg ctl_reg_gp_hilo_pla23pla16M2T2_4;
reg ctl_reg_gp_sel_pla23pla16M2T3_5;
reg ctl_reg_gp_hilo_pla23pla16M2T3_6;
reg ctl_reg_gp_sel_pla23pla16M3T1_5;
reg ctl_reg_gp_hilo_pla23pla16M3T1_6;
reg ctl_reg_gp_sel_pla23pla16M3T2_3;
reg ctl_reg_gp_hilo_pla23pla16M3T2_4;
reg ctl_reg_gp_sel_pla23npla16M2T1_3;
reg ctl_reg_gp_hilo_pla23npla16M2T1_4;
reg ctl_reg_gp_sel_pla23npla16M2T2_3;
reg ctl_reg_gp_hilo_pla23npla16M2T2_4;
reg ctl_reg_gp_sel_pla23npla16M2T3_5;
reg ctl_reg_gp_hilo_pla23npla16M2T3_6;
reg ctl_reg_gp_sel_pla23npla16M3T1_3;
reg ctl_reg_gp_hilo_pla23npla16M3T1_4;
reg ctl_reg_gp_sel_pla23npla16M3T2_3;
reg ctl_reg_gp_hilo_pla23npla16M3T2_4;
reg ctl_reg_gp_sel_pla23npla16M3T3_4;
reg ctl_reg_gp_hilo_pla23npla16M3T3_5;
reg ctl_reg_gp_sel_pla10M2T1_3;
reg ctl_reg_gp_hilo_pla10M2T1_4;
reg ctl_reg_gp_sel_pla10M2T2_3;
reg ctl_reg_gp_hilo_pla10M2T2_4;
reg ctl_reg_sys_hilo_pla10M2T3_6;
reg ctl_reg_gp_sel_pla10M3T1_3;
reg ctl_reg_gp_hilo_pla10M3T1_4;
reg ctl_reg_gp_sel_pla10M3T2_3;
reg ctl_reg_gp_hilo_pla10M3T2_4;
reg ctl_reg_sys_hilo_pla10M3T3_4;
reg ctl_reg_gp_sel_pla10M3T4_4;
reg ctl_reg_gp_hilo_pla10M3T4_5;
reg ctl_reg_gp_sel_pla10M4T1_5;
reg ctl_reg_gp_hilo_pla10M4T1_6;
reg ctl_reg_gp_sel_pla10M4T2_3;
reg ctl_reg_gp_hilo_pla10M4T2_4;
reg ctl_reg_gp_sel_pla10M4T3_5;
reg ctl_reg_gp_hilo_pla10M4T3_6;
reg ctl_reg_gp_sel_pla10M5T1_5;
reg ctl_reg_gp_hilo_pla10M5T1_6;
reg ctl_reg_gp_sel_pla10M5T2_3;
reg ctl_reg_gp_hilo_pla10M5T2_4;
reg ctl_reg_sys_hilo_pla10M5T3_3;
reg ctl_reg_gp_sel_pla10M5T4_2;
reg ctl_reg_gp_hilo_pla10M5T4_3;
reg ctl_pf_sel_pla12M1T1_12;
reg ctl_reg_gp_sel_pla12M1T2_2;
reg ctl_reg_gp_hilo_pla12M1T2_3;
reg ctl_reg_gp_sel_pla12M1T3_1;
reg ctl_reg_gp_hilo_pla12M1T3_2;
reg ctl_reg_gp_sel_pla12M2T1_2;
reg ctl_reg_gp_hilo_pla12M2T1_3;
reg ctl_reg_gp_sel_pla12M2T2_3;
reg ctl_reg_gp_hilo_pla12M2T2_4;
reg ctl_reg_gp_sel_pla12M3T1_2;
reg ctl_reg_gp_hilo_pla12M3T1_3;
reg ctl_reg_gp_sel_pla12M3T2_3;
reg ctl_reg_gp_hilo_pla12M3T2_4;
reg ctl_reg_gp_sel_pla12M3T3_2;
reg ctl_reg_gp_hilo_pla12M3T3_3;
reg ctl_reg_gp_sel_pla12M3T4_2;
reg ctl_reg_gp_hilo_pla12M3T4_3;
reg ctl_reg_sys_hilo_pla12M4T1_2;
reg ctl_reg_sys_hilo_pla12M4T2_3;
reg ctl_reg_sys_hilo_pla12M4T3_2;
reg ctl_reg_sys_hilo_pla12M4T4_3;
reg ctl_pf_sel_pla11M1T1_11;
reg ctl_reg_gp_sel_pla11M1T2_2;
reg ctl_reg_gp_hilo_pla11M1T2_3;
reg ctl_reg_gp_sel_pla11M1T3_1;
reg ctl_reg_gp_hilo_pla11M1T3_2;
reg ctl_reg_gp_sel_pla11M2T1_2;
reg ctl_reg_gp_hilo_pla11M2T1_3;
reg ctl_reg_gp_sel_pla11M2T2_3;
reg ctl_reg_gp_hilo_pla11M2T2_4;
reg ctl_reg_gp_sel_pla11M3T3_1;
reg ctl_reg_gp_hilo_pla11M3T3_2;
reg ctl_reg_gp_sel_pla11M3T4_2;
reg ctl_reg_gp_hilo_pla11M3T4_3;
reg ctl_reg_sys_hilo_pla11M4T1_2;
reg ctl_reg_sys_hilo_pla11M4T2_3;
reg ctl_reg_sys_hilo_pla11M4T3_2;
reg ctl_reg_sys_hilo_pla11M4T4_3;
reg ctl_reg_gp_sel_pla65npla52M1T2_2;
reg ctl_reg_gp_hilo_pla65npla52M1T2_3;
reg ctl_reg_gp_sel_pla65npla52M1T3_1;
reg ctl_reg_gp_hilo_pla65npla52M1T3_2;
reg ctl_reg_gp_sel_pla65npla52M1T4_3;
reg ctl_reg_gp_hilo_pla65npla52M1T4_4;
reg ctl_reg_gp_sel_pla64M1T2_2;
reg ctl_reg_gp_hilo_pla64M1T2_3;
reg ctl_reg_gp_sel_pla64M1T3_1;
reg ctl_reg_gp_hilo_pla64M1T3_2;
reg ctl_reg_gp_sel_pla64M1T4_4;
reg ctl_reg_gp_hilo_pla64M1T4_5;
reg ctl_reg_sys_hilo_pla64M2T1_3;
reg ctl_reg_sys_hilo_pla64M2T2_4;
reg ctl_reg_gp_sel_use_ixiypla52M1T3_1;
reg ctl_reg_gp_hilo_use_ixiypla52M1T3_2;
reg ctl_reg_sys_hilo_use_ixiypla52M2T1_3;
reg ctl_reg_sys_hilo_use_ixiypla52M2T2_4;
reg ctl_reg_gp_sel_nuse_ixiypla52M1T2_2;
reg ctl_reg_gp_hilo_nuse_ixiypla52M1T2_3;
reg ctl_reg_gp_sel_nuse_ixiypla52M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla52M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla52M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla52M2T1_3;
reg ctl_reg_sys_hilo_nuse_ixiypla52M2T2_4;
reg ctl_reg_gp_sel_nuse_ixiypla52M4T2_2;
reg ctl_reg_gp_hilo_nuse_ixiypla52M4T2_3;
reg ctl_reg_gp_sel_pla66npla53M1T1_2;
reg ctl_reg_gp_hilo_pla66npla53M1T1_3;
reg ctl_pf_sel_pla66npla53M1T1_15;
reg ctl_reg_gp_sel_pla66npla53M1T2_2;
reg ctl_reg_gp_hilo_pla66npla53M1T2_3;
reg ctl_reg_gp_sel_pla66npla53M1T3_1;
reg ctl_reg_gp_hilo_pla66npla53M1T3_2;
reg ctl_reg_gp_sel_pla66npla53M1T4nop4op5nop3_1;
reg ctl_reg_gp_hilo_pla66npla53M1T4nop4op5nop3_2;
reg ctl_reg_gp_sel_use_ixiypla53M1T3_1;
reg ctl_reg_gp_hilo_use_ixiypla53M1T3_2;
reg ctl_reg_sys_hilo_use_ixiypla53M2T1_3;
reg ctl_reg_sys_hilo_use_ixiypla53M2T2_4;
reg ctl_reg_gp_sel_nuse_ixiypla53M1T2_2;
reg ctl_reg_gp_hilo_nuse_ixiypla53M1T2_3;
reg ctl_reg_gp_sel_nuse_ixiypla53M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla53M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla53M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla53M2T1_3;
reg ctl_pf_sel_nuse_ixiypla53M2T4_14;
reg ctl_pf_sel_nuse_ixiypla53M4T4_14;
reg ctl_reg_gp_sel_pla69M1T2_2;
reg ctl_reg_gp_hilo_pla69M1T2_3;
reg ctl_reg_gp_sel_pla69M1T3_1;
reg ctl_reg_gp_hilo_pla69M1T3_2;
reg ctl_reg_gp_sel_pla69M1T4_3;
reg ctl_reg_gp_hilo_pla69M1T4_4;
reg ctl_reg_gp_sel_pla69M2T1_1;
reg ctl_reg_gp_hilo_pla69M2T1_2;
reg ctl_reg_sys_hilo_pla69M2T2_3;
reg ctl_reg_gp_sel_pla69M2T3_1;
reg ctl_reg_gp_hilo_pla69M2T3_2;
reg ctl_reg_gp_sel_pla69M2T4_2;
reg ctl_reg_gp_hilo_pla69M2T4_3;
reg ctl_reg_sys_hilo_pla69M3T1_2;
reg ctl_reg_sys_hilo_pla69M3T1_7;
reg ctl_reg_gp_sel_pla69M3T2_2;
reg ctl_reg_gp_hilo_pla69M3T2_3;
reg ctl_reg_gp_sel_op3pla68M1T2_2;
reg ctl_reg_gp_hilo_op3pla68M1T2_3;
reg ctl_reg_gp_sel_op3pla68M1T3_1;
reg ctl_reg_gp_hilo_op3pla68M1T3_2;
reg ctl_reg_gp_sel_op3pla68M1T4_3;
reg ctl_reg_gp_hilo_op3pla68M1T4_4;
reg ctl_reg_gp_sel_op3pla68M2T1_1;
reg ctl_reg_gp_hilo_op3pla68M2T1_2;
reg ctl_reg_sys_hilo_op3pla68M2T2_3;
reg ctl_reg_gp_sel_op3pla68M2T3_1;
reg ctl_reg_gp_hilo_op3pla68M2T3_2;
reg ctl_reg_gp_sel_op3pla68M2T4_2;
reg ctl_reg_gp_hilo_op3pla68M2T4_3;
reg ctl_reg_sys_hilo_op3pla68M3T1_2;
reg ctl_reg_sys_hilo_op3pla68M3T1_7;
reg ctl_pf_sel_op3pla68M3T1_18;
reg ctl_reg_gp_sel_op3pla68M3T2_2;
reg ctl_reg_gp_hilo_op3pla68M3T2_3;
reg ctl_reg_gp_sel_nop3pla68M1T2_2;
reg ctl_reg_gp_hilo_nop3pla68M1T2_3;
reg ctl_reg_gp_sel_nop3pla68M1T3_1;
reg ctl_reg_gp_hilo_nop3pla68M1T3_2;
reg ctl_reg_gp_sel_nop3pla68M1T4_3;
reg ctl_reg_gp_hilo_nop3pla68M1T4_4;
reg ctl_reg_gp_sel_nop3pla68M2T1_1;
reg ctl_reg_gp_hilo_nop3pla68M2T1_2;
reg ctl_reg_sys_hilo_nop3pla68M2T2_3;
reg ctl_reg_gp_sel_nop3pla68M2T3_1;
reg ctl_reg_gp_hilo_nop3pla68M2T3_2;
reg ctl_reg_gp_sel_nop3pla68M2T4_2;
reg ctl_reg_gp_hilo_nop3pla68M2T4_3;
reg ctl_reg_sys_hilo_nop3pla68M3T1_2;
reg ctl_reg_sys_hilo_nop3pla68M3T1_7;
reg ctl_pf_sel_nop3pla68M3T1_20;
reg ctl_reg_gp_sel_nop3pla68M3T2_2;
reg ctl_reg_gp_hilo_nop3pla68M3T2_3;
reg ctl_reg_gp_sel_pla9M1T4_2;
reg ctl_reg_gp_hilo_pla9M1T4_3;
reg ctl_reg_gp_sel_pla9M1T5_2;
reg ctl_reg_gp_hilo_pla9M1T5_3;
reg ctl_reg_gp_sel_pla77M1T1_2;
reg ctl_reg_gp_hilo_pla77M1T1_3;
reg ctl_pf_sel_pla77M1T1_14;
reg ctl_reg_gp_sel_pla77M1T2_2;
reg ctl_reg_gp_hilo_pla77M1T2_3;
reg ctl_reg_gp_sel_pla77M1T3_1;
reg ctl_reg_gp_hilo_pla77M1T3_2;
reg ctl_reg_gp_sel_pla81M1T1_2;
reg ctl_reg_gp_hilo_pla81M1T1_3;
reg ctl_reg_gp_sel_pla81M1T2_2;
reg ctl_reg_gp_hilo_pla81M1T2_3;
reg ctl_reg_gp_sel_pla81M1T3_1;
reg ctl_reg_gp_hilo_pla81M1T3_2;
reg ctl_reg_gp_sel_pla82M1T1_2;
reg ctl_reg_gp_hilo_pla82M1T1_3;
reg ctl_pf_sel_pla82M1T1_16;
reg ctl_reg_gp_sel_pla82M1T2_2;
reg ctl_reg_gp_hilo_pla82M1T2_3;
reg ctl_reg_gp_sel_pla82M1T3_1;
reg ctl_reg_gp_hilo_pla82M1T3_2;
reg ctl_reg_gp_sel_pla89M1T2_2;
reg ctl_reg_gp_hilo_pla89M1T2_3;
reg ctl_reg_gp_sel_pla89M1T3_1;
reg ctl_reg_gp_hilo_pla89M1T3_2;
reg ctl_reg_gp_sel_pla92M1T2_2;
reg ctl_reg_gp_hilo_pla92M1T2_3;
reg ctl_reg_gp_sel_pla92M1T3_1;
reg ctl_reg_gp_hilo_pla92M1T3_2;
reg ctl_reg_gp_sel_pla25M1T1_2;
reg ctl_reg_gp_hilo_pla25M1T1_3;
reg ctl_reg_gp_sel_pla25M1T2_2;
reg ctl_reg_gp_hilo_pla25M1T2_3;
reg ctl_reg_gp_sel_pla25M1T3_1;
reg ctl_reg_gp_hilo_pla25M1T3_2;
reg ctl_reg_gp_sel_pla25M1T4_3;
reg ctl_reg_gp_hilo_pla25M1T4_4;
reg ctl_reg_gp_sel_nuse_ixiypla70npla55M1T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T1_3;
reg ctl_pf_sel_nuse_ixiypla70npla55M1T1_20;
reg ctl_reg_gp_sel_nuse_ixiypla70npla55M1T2_2;
reg ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T2_3;
reg ctl_reg_gp_sel_nuse_ixiypla70npla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla70npla55M1T4_3;
reg ctl_reg_gp_hilo_nuse_ixiypla70npla55M1T4_4;
reg ctl_reg_sys_hilo_nuse_ixiypla70npla55M4T1_3;
reg ctl_pf_sel_nuse_ixiypla70npla55M5T1_19;
reg ctl_reg_gp_sel_nuse_ixiypla70pla55M1T2_2;
reg ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T2_3;
reg ctl_reg_gp_sel_nuse_ixiypla70pla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla70pla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla70pla55M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla70pla55M2T1_3;
reg ctl_pf_sel_nuse_ixiypla70pla55M3T1_19;
reg ctl_reg_sys_hilo_nuse_ixiypla70pla55M4T1_3;
reg ctl_pf_sel_nuse_ixiypla70pla55M5T1_19;
reg ctl_reg_gp_sel_pla15op3M1T1_2;
reg ctl_reg_gp_hilo_pla15op3M1T1_3;
reg ctl_pf_sel_pla15op3M1T1_18;
reg ctl_reg_gp_sel_pla15op3M1T2_2;
reg ctl_reg_gp_hilo_pla15op3M1T2_3;
reg ctl_reg_gp_sel_pla15op3M1T3_1;
reg ctl_reg_gp_hilo_pla15op3M1T3_2;
reg ctl_reg_gp_sel_pla15op3M2T1_2;
reg ctl_reg_gp_hilo_pla15op3M2T1_3;
reg ctl_reg_sys_hilo_pla15op3M2T2_4;
reg ctl_reg_gp_sel_pla15nop3M1T1_2;
reg ctl_reg_gp_hilo_pla15nop3M1T1_3;
reg ctl_pf_sel_pla15nop3M1T1_18;
reg ctl_reg_gp_sel_pla15nop3M1T2_2;
reg ctl_reg_gp_hilo_pla15nop3M1T2_3;
reg ctl_reg_gp_sel_pla15nop3M1T3_1;
reg ctl_reg_gp_hilo_pla15nop3M1T3_2;
reg ctl_reg_gp_sel_pla15nop3M2T1_2;
reg ctl_reg_gp_hilo_pla15nop3M2T1_3;
reg ctl_reg_sys_hilo_pla15nop3M2T2_4;
reg ctl_reg_gp_sel_pla15nop3M3T3_1;
reg ctl_reg_gp_hilo_pla15nop3M3T3_2;
reg ctl_pf_sel_nuse_ixiypla72npla55M1T1_10;
reg ctl_reg_gp_sel_nuse_ixiypla72npla55M1T2_2;
reg ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T2_3;
reg ctl_reg_gp_sel_nuse_ixiypla72npla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla72npla55M1T4_3;
reg ctl_reg_gp_hilo_nuse_ixiypla72npla55M1T4_4;
reg ctl_pf_sel_nuse_ixiypla72pla55M1T1_10;
reg ctl_reg_gp_sel_nuse_ixiypla72pla55M1T2_2;
reg ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T2_3;
reg ctl_reg_gp_sel_nuse_ixiypla72pla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla72pla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla72pla55M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla72pla55M2T1_3;
reg ctl_reg_sys_hilo_nuse_ixiypla72pla55M2T3_3;
reg ctl_reg_sys_hilo_nuse_ixiypla72pla55M4T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla74npla55M1T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla74npla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla74npla55M1T4_3;
reg ctl_reg_gp_hilo_nuse_ixiypla74npla55M1T4_4;
reg ctl_reg_sys_hilo_nuse_ixiypla74npla55M4T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla74pla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla74pla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla74pla55M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla74pla55M2T1_3;
reg ctl_reg_sys_hilo_nuse_ixiypla74pla55M4T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla73npla55M1T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla73npla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla73npla55M1T4_3;
reg ctl_reg_gp_hilo_nuse_ixiypla73npla55M1T4_4;
reg ctl_reg_sys_hilo_nuse_ixiypla73npla55M4T1_3;
reg ctl_reg_gp_sel_nuse_ixiypla73pla55M1T3_1;
reg ctl_reg_gp_hilo_nuse_ixiypla73pla55M1T3_2;
reg ctl_reg_gp_sel_nuse_ixiypla73pla55M2T1_2;
reg ctl_reg_gp_hilo_nuse_ixiypla73pla55M2T1_3;
reg ctl_reg_sys_hilo_nuse_ixiypla73pla55M4T1_3;
reg ctl_reg_gp_sel_pla37npla28M1T1_2;
reg ctl_reg_gp_hilo_pla37npla28M1T1_3;
reg ctl_reg_sys_hilo_pla37npla28M2T1_3;
reg ctl_reg_sys_hilo_pla37npla28M2T2_4;
reg ctl_reg_gp_sel_pla37npla28M3T1_2;
reg ctl_reg_gp_hilo_pla37npla28M3T1_3;
reg ctl_reg_gp_sel_pla27npla34M1T1_2;
reg ctl_reg_gp_hilo_pla27npla34M1T1_3;
reg ctl_pf_sel_pla27npla34M1T1_20;
reg ctl_reg_gp_sel_pla27npla34M1T2_2;
reg ctl_reg_gp_hilo_pla27npla34M1T2_3;
reg ctl_reg_gp_sel_pla27npla34M1T3_1;
reg ctl_reg_gp_hilo_pla27npla34M1T3_2;
reg ctl_reg_gp_sel_pla27npla34M2T1_2;
reg ctl_reg_gp_hilo_pla27npla34M2T1_3;
reg ctl_reg_sys_hilo_pla37pla28M2T1_3;
reg ctl_reg_sys_hilo_pla37pla28M2T2_4;
reg ctl_reg_gp_sel_pla37pla28M2T3_4;
reg ctl_reg_gp_hilo_pla37pla28M2T3_5;
reg ctl_reg_gp_sel_pla37pla28M3T1_3;
reg ctl_reg_gp_hilo_pla37pla28M3T1_4;
reg ctl_reg_gp_sel_pla27pla34M1T4nop4op5nop3_1;
reg ctl_reg_gp_hilo_pla27pla34M1T4nop4op5nop3_2;
reg ctl_reg_gp_sel_pla27pla34M2T1_2;
reg ctl_reg_gp_hilo_pla27pla34M2T1_3;
reg ctl_pf_sel_pla91pla21M1T1_8;
reg ctl_reg_gp_sel_pla91pla21M1T2_2;
reg ctl_reg_gp_hilo_pla91pla21M1T2_3;
reg ctl_reg_gp_sel_pla91pla21M1T3_1;
reg ctl_reg_gp_hilo_pla91pla21M1T3_2;
reg ctl_reg_gp_sel_pla91pla21M2T1_2;
reg ctl_reg_gp_hilo_pla91pla21M2T1_3;
reg ctl_reg_gp_sel_pla91pla21M2T2_2;
reg ctl_reg_gp_hilo_pla91pla21M2T2_3;
reg ctl_reg_gp_sel_pla91pla21M2T3_3;
reg ctl_reg_gp_hilo_pla91pla21M2T3_4;
reg ctl_reg_gp_sel_pla91pla21M3T1_2;
reg ctl_reg_gp_hilo_pla91pla21M3T1_3;
reg ctl_reg_gp_sel_pla91pla21M3T2_3;
reg ctl_reg_gp_hilo_pla91pla21M3T2_4;
reg ctl_reg_sys_hilo_pla91pla21M4T1_2;
reg ctl_reg_sys_hilo_pla91pla21M4T2_3;
reg ctl_reg_sys_hilo_pla91pla21M4T3_2;
reg ctl_reg_sys_hilo_pla91pla21M4T4_3;
reg ctl_pf_sel_pla91pla20M1T1_9;
reg ctl_reg_gp_sel_pla91pla20M1T2_2;
reg ctl_reg_gp_hilo_pla91pla20M1T2_3;
reg ctl_reg_gp_sel_pla91pla20M1T3_1;
reg ctl_reg_gp_hilo_pla91pla20M1T3_2;
reg ctl_reg_gp_sel_pla91pla20M1T4_2;
reg ctl_reg_gp_hilo_pla91pla20M1T4_3;
reg ctl_reg_gp_sel_pla91pla20M1T5_4;
reg ctl_reg_gp_hilo_pla91pla20M1T5_5;
reg ctl_reg_gp_sel_pla91pla20M2T1_2;
reg ctl_reg_gp_hilo_pla91pla20M2T1_3;
reg ctl_reg_gp_sel_pla91pla20M2T2_3;
reg ctl_reg_gp_hilo_pla91pla20M2T2_4;
reg ctl_reg_gp_sel_pla91pla20M2T3_4;
reg ctl_reg_gp_hilo_pla91pla20M2T3_5;
reg ctl_reg_gp_sel_pla91pla20M3T1_2;
reg ctl_reg_gp_hilo_pla91pla20M3T1_3;
reg ctl_reg_sys_hilo_pla91pla20M4T1_2;
reg ctl_reg_sys_hilo_pla91pla20M4T2_3;
reg ctl_reg_sys_hilo_pla91pla20M4T3_2;
reg ctl_reg_sys_hilo_pla91pla20M4T4_3;
reg ctl_reg_sys_hilo_pla29M2T1_3;
reg ctl_reg_sys_hilo_pla29M2T2_4;
reg ctl_reg_sys_hilo_pla29M2T3_6;
reg ctl_reg_sys_hilo_pla29M3T1_3;
reg ctl_reg_sys_hilo_pla29M3T2_4;
reg ctl_reg_sys_hilo_pla29M3T3_4;
reg ctl_reg_sys_hilo_pla29M3T3_9;
reg ctl_reg_gp_sel_pla43M1T3_1;
reg ctl_reg_gp_hilo_pla43M1T3_2;
reg ctl_reg_sys_hilo_pla43M2T1_3;
reg ctl_reg_sys_hilo_pla43M2T2_4;
reg ctl_reg_sys_hilo_pla43M2T3_6;
reg ctl_reg_sys_hilo_pla43M3T1_3;
reg ctl_reg_sys_hilo_pla43M3T2_4;
reg ctl_reg_sys_hilo_pla43M3T3_5;
reg ctl_reg_sys_hilo_pla43M3T3_10;
reg ctl_reg_gp_sel_pla47M1T3_1;
reg ctl_reg_gp_hilo_pla47M1T3_2;
reg ctl_reg_sys_hilo_pla47M2T1_3;
reg ctl_reg_sys_hilo_pla47M2T2_4;
reg ctl_reg_sys_hilo_pla47M3T2_2;
reg ctl_reg_sys_hilo_pla47M3T3_3;
reg ctl_reg_sys_hilo_pla47M3T4_2;
reg ctl_reg_sys_hilo_pla47M3T5_3;
reg ctl_reg_sys_hilo_pla47M3T5_8;
reg ctl_reg_gp_sel_pla48M1T3_1;
reg ctl_reg_gp_hilo_pla48M1T3_2;
reg ctl_reg_sys_hilo_pla48M2T1_3;
reg ctl_reg_sys_hilo_pla48M2T2_4;
reg ctl_reg_sys_hilo_pla48M3T2_2;
reg ctl_reg_sys_hilo_pla48M3T3_3;
reg ctl_reg_sys_hilo_pla48M3T4_2;
reg ctl_reg_sys_hilo_pla48M3T5_3;
reg ctl_reg_sys_hilo_pla48M3T5_8;
reg ctl_reg_gp_sel_pla6M1T4_3;
reg ctl_reg_gp_hilo_pla6M1T4_4;
reg ctl_reg_gp_sel_pla26M1T3_1;
reg ctl_reg_gp_hilo_pla26M1T3_2;
reg ctl_reg_gp_sel_pla26M1T4_2;
reg ctl_reg_gp_hilo_pla26M1T4_3;
reg ctl_reg_gp_sel_pla26M1T5_4;
reg ctl_reg_gp_hilo_pla26M1T5_5;
reg ctl_reg_sys_hilo_pla26M2T1_3;
reg ctl_reg_sys_hilo_pla26M2T2_4;
reg ctl_reg_sys_hilo_pla26M3T2_2;
reg ctl_reg_sys_hilo_pla26M3T3_3;
reg ctl_reg_sys_hilo_pla26M3T4_2;
reg ctl_reg_sys_hilo_pla26M3T5_3;
reg ctl_reg_sys_hilo_pla26M3T5_8;
reg ctl_reg_sys_hilo_pla24M2T1_3;
reg ctl_reg_sys_hilo_pla24M2T2_4;
reg ctl_reg_sys_hilo_pla24M2T3_6;
reg ctl_reg_sys_hilo_pla24M3T1_3;
reg ctl_reg_sys_hilo_pla24M3T2_4;
reg ctl_reg_sys_hilo_pla24M3T3_4;
reg ctl_reg_gp_sel_pla24M3T4_4;
reg ctl_reg_gp_hilo_pla24M3T4_5;
reg ctl_reg_sys_hilo_pla24M4T1_6;
reg ctl_reg_gp_sel_pla24M4T2_3;
reg ctl_reg_gp_hilo_pla24M4T2_4;
reg ctl_reg_gp_sel_pla24M4T3_5;
reg ctl_reg_gp_hilo_pla24M4T3_6;
reg ctl_reg_sys_hilo_pla24M5T1_6;
reg ctl_reg_gp_sel_pla24M5T2_3;
reg ctl_reg_gp_hilo_pla24M5T2_4;
reg ctl_reg_sys_hilo_pla24M5T3_4;
reg ctl_reg_gp_sel_pla42M1T3_1;
reg ctl_reg_gp_hilo_pla42M1T3_2;
reg ctl_reg_sys_hilo_pla42M2T1_3;
reg ctl_reg_sys_hilo_pla42M2T2_4;
reg ctl_reg_sys_hilo_pla42M2T3_6;
reg ctl_reg_sys_hilo_pla42M3T1_3;
reg ctl_reg_sys_hilo_pla42M3T2_4;
reg ctl_reg_sys_hilo_pla42M3T3_6;
reg ctl_reg_gp_sel_pla42M3T4_4;
reg ctl_reg_gp_hilo_pla42M3T4_5;
reg ctl_reg_sys_hilo_pla42M4T1_6;
reg ctl_reg_gp_sel_pla42M4T2_3;
reg ctl_reg_gp_hilo_pla42M4T2_4;
reg ctl_reg_gp_sel_pla42M4T3_5;
reg ctl_reg_gp_hilo_pla42M4T3_6;
reg ctl_reg_sys_hilo_pla42M5T1_6;
reg ctl_reg_gp_sel_pla42M5T2_3;
reg ctl_reg_gp_hilo_pla42M5T2_4;
reg ctl_reg_sys_hilo_pla42M5T3_4;
reg ctl_reg_gp_sel_pla35M2T1_3;
reg ctl_reg_gp_hilo_pla35M2T1_4;
reg ctl_reg_gp_sel_pla35M2T2_3;
reg ctl_reg_gp_hilo_pla35M2T2_4;
reg ctl_reg_sys_hilo_pla35M2T3_6;
reg ctl_reg_gp_sel_pla35M3T1_3;
reg ctl_reg_gp_hilo_pla35M3T1_4;
reg ctl_reg_gp_sel_pla35M3T2_3;
reg ctl_reg_gp_hilo_pla35M3T2_4;
reg ctl_reg_sys_hilo_pla35M3T3_4;
reg ctl_reg_sys_hilo_pla35M3T3_9;
reg ctl_reg_gp_sel_pla45M1T3_1;
reg ctl_reg_gp_hilo_pla45M1T3_2;
reg ctl_reg_gp_sel_pla45M2T1_3;
reg ctl_reg_gp_hilo_pla45M2T1_4;
reg ctl_reg_gp_sel_pla45M2T2_3;
reg ctl_reg_gp_hilo_pla45M2T2_4;
reg ctl_reg_sys_hilo_pla45M2T3_6;
reg ctl_reg_gp_sel_pla45M3T1_3;
reg ctl_reg_gp_hilo_pla45M3T1_4;
reg ctl_reg_gp_sel_pla45M3T2_3;
reg ctl_reg_gp_hilo_pla45M3T2_4;
reg ctl_reg_sys_hilo_pla45M3T3_4;
reg ctl_reg_sys_hilo_pla45M3T3_9;
reg ctl_reg_gp_sel_pla46M2T1_3;
reg ctl_reg_gp_hilo_pla46M2T1_4;
reg ctl_reg_gp_sel_pla46M2T2_3;
reg ctl_reg_gp_hilo_pla46M2T2_4;
reg ctl_reg_sys_hilo_pla46M2T3_6;
reg ctl_reg_gp_sel_pla46M3T1_3;
reg ctl_reg_gp_hilo_pla46M3T1_4;
reg ctl_reg_gp_sel_pla46M3T2_3;
reg ctl_reg_gp_hilo_pla46M3T2_4;
reg ctl_reg_sys_hilo_pla46M3T3_4;
reg ctl_reg_sys_hilo_pla46M3T3_9;
reg ctl_reg_sys_hilo_pla56M1T3_3;
reg ctl_reg_gp_sel_pla56M1T5_4;
reg ctl_reg_gp_hilo_pla56M1T5_5;
reg ctl_reg_sys_hilo_pla56M2T1_6;
reg ctl_reg_gp_sel_pla56M2T2_3;
reg ctl_reg_gp_hilo_pla56M2T2_4;
reg ctl_reg_gp_sel_pla56M2T3_5;
reg ctl_reg_gp_hilo_pla56M2T3_6;
reg ctl_reg_sys_hilo_pla56M3T1_6;
reg ctl_reg_gp_sel_pla56M3T2_3;
reg ctl_reg_gp_hilo_pla56M3T2_4;
reg ctl_reg_sys_hilo_pla56M3T3_6;
reg ctl_reg_sys_hilo_pla56M4T1_3;
reg ctl_reg_sys_hilo_pla56M4T3_6;
reg ctl_reg_sys_hilo_pla56M5T1_3;
reg ctl_reg_sys_hilo_pla56M5T3_4;
reg ctl_reg_sys_hilo_pla56M5T3_9;
reg ctl_reg_gp_sel_pla49M1T3_1;
reg ctl_reg_gp_hilo_pla49M1T3_2;
reg ctl_reg_sys_hilo_pla49M2T1_3;
reg ctl_reg_sys_hilo_pla49M2T2_4;
reg ctl_reg_sys_hilo_pla49M3T1_3;
reg ctl_reg_sys_hilo_pla49M3T2_4;
reg ctl_pf_sel_pla76M1T1_2;
reg ctl_reg_gp_sel_pla78M1T1_2;
reg ctl_reg_gp_hilo_pla78M1T1_3;
reg ctl_pf_sel_pla78M1T1_8;
reg ctl_reg_gp_sel_pla79M1T1_2;
reg ctl_reg_gp_hilo_pla79M1T1_3;
reg ctl_pf_sel_pla79M1T1_8;
reg ctl_reg_gp_sel_pla80M1T1_2;
reg ctl_reg_gp_hilo_pla80M1T1_3;
reg ctl_pf_sel_pla80M1T1_8;
reg ctl_reg_gp_sel_pla84M1T1_2;
reg ctl_reg_gp_hilo_pla84M1T1_3;
reg ctl_pf_sel_pla84M1T1_8;
reg ctl_reg_gp_sel_pla85M1T1_2;
reg ctl_reg_gp_hilo_pla85M1T1_3;
reg ctl_pf_sel_pla85M1T1_8;
reg ctl_reg_gp_sel_pla86M1T1_2;
reg ctl_reg_gp_hilo_pla86M1T1_3;
reg ctl_pf_sel_pla86M1T1_8;
reg ctl_reg_gp_sel_pla88M1T1_2;
reg ctl_reg_gp_hilo_pla88M1T1_3;
reg ctl_pf_sel_pla88M1T1_8;
reg ctl_reg_gp_sel_ixy_dT2_1;
reg ctl_reg_gp_hilo_ixy_dT2_2;
reg ctl_reg_sys_hilo_ixy_dT3_3;
reg ctl_reg_gp_sel_ixy_dT4_1;
reg ctl_reg_gp_hilo_ixy_dT4_2;
reg ctl_reg_sys_hilo_ixy_dT5_2;
reg ctl_reg_sys_hilo_ixy_dT5_7;
reg ctl_reg_sys_hilo_1M1T1_3;
reg ctl_reg_sys_hilo_1M1T2_2;
reg ctl_reg_sys_hilo_1M1T3_3;
reg ctl_reg_sys_hilo_setM1_2;
